���*      }�(K�nicobar�K�north and middle andaman�K�south andaman�K	�	anantapur�K
�chittoor�K�east godavari�K�guntur�K�krishna�K�kurnool�K�prakasam�K�sri potti sriramulu nellore�K�
srikakulam�K�visakhapatnam�K�vizianagaram�K�west godavari�K�ysr district, kadapa (cuddapah)�K�anjaw�K�	changlang�K�dibang valley�K�east kameng�K*�
east siang�K�itanagar capital complex�K�kamle�K�	kra daadi�K�kurung kumey�K!�	lepa rada�K�lohit�K(�longding�K�lower dibang valley�K�lower siang�K �lower subansiri�K$�namsai�K�pakke kessang�K'�
papum pare�K#�shi yomi�K%�siang�K�tawang�K�tirap�K"�upper siang�K)�upper subansiri�K�west kameng�K&�
west siang�K.�baksa�K/�barpeta�M��	biswanath�K9�
bongaigaon�KB�cachar�M��	charaideo�K:�chirang�K0�darrang�K>�dhemaji�K;�dhubri�K+�	dibrugarh�KC�
dima hasao�K<�goalpara�K5�golaghat�KD�
hailakandi�M��hojai�K6�jorhat�K1�kamrup metropolitan�K2�kamrup rural�K3�karbi-anglong�KE�	karimganj�K=�	kokrajhar�K?�	lakhimpur�M��majuli�K7�morigaon�K8�nagaon�K4�nalbari�K,�	sivasagar�K@�sonitpur�M �south salmara mankachar�K-�tinsukia�KA�udalguri�M�west karbi anglong�KJ�araria�KN�arwal�KM�
aurangabad�KS�banka�Kb�	begusarai�KR�	bhagalpur�Kc�bhojpur�Kd�buxar�K^�	darbhanga�Ki�east champaran�KO�gaya�Kh�	gopalganj�Kk�jamui�K[�	jehanabad�KP�kaimur�KK�katihar�Ke�khagaria�KL�
kishanganj�KT�
lakhisarai�KF�	madhepura�K_�	madhubani�KU�munger�KV�muzaffarpur�KZ�nalanda�K\�nawada�Ka�patna�KI�purnia�KQ�rohtas�KG�saharsa�K`�
samastipur�Kf�saran�K]�
sheikhpura�KW�sheohar�KX�	sitamarhi�Kg�siwan�KH�supaul�KY�vaishali�Kj�west champaran�Kl�
chandigarh�Kn�balod�Ko�baloda bazar�Kp�	balrampur�Kq�bastar�Kr�bemetara�Ks�bijapur�Kt�bilaspur�Ku�	dantewada�Kv�dhamtari�Kw�durg�Kx�	gariaband�K��gaurela pendra marwahi �Ky�janjgir-champa�Kz�jashpur�K{�kanker�K��kawardha�K|�	kondagaon�K}�korba�K~�koriya�K�
mahasamund�K��mungeli�K��
narayanpur�K��raigarh�Km�raipur�K��rajnandgaon�K��sukma�K��surajpur�K��surguja�K��dadra and nagar haveli�K��daman�K��diu�K��central delhi�K��
east delhi�K��	new delhi�K��north delhi�K��north east delhi�K��north west delhi�K��shahdara�K��south delhi�K��south east delhi�K��south west delhi�K��
west delhi�K��	north goa�K��	south goa�K��	ahmedabad�M�ahmedabad corporation�K��amreli�K��anand�K��aravalli�K��banaskantha�K��bharuch�K��	bhavnagar�M�bhavnagar corporation�K��botad�K��chhotaudepur�K��dahod�K��dang�K��devbhumi dwaraka�K��gandhinagar�M�gandhinagar corporation�K��gir somnath�K��jamnagar�M�jamnagar corporation�K��junagadh�M�junagadh corporation�K��kheda�K��kutch�K��	mahisagar�K��mehsana�K��morbi�K��narmada�K��navsari�K��
panchmahal�K��patan�K��	porbandar�K��rajkot�M�rajkot corporation�K��sabarkantha�K��surat�M�surat corporation�K��surendranagar�K��tapi�K��vadodara�M	�vadodara corporation�K��valsad�K��ambala�KȌbhiwani�KɌcharkhi dadri�Kǌ	faridabad�KČ	fatehabad�K��gurgaon�K��hisar�K��jhajjar�Ǩjind�K��kaithal�Kˌkarnal�K��kurukshetra�KΌmahendragarh�K͌nuh�Kόpalwal�K��	panchkula�KÌpanipat�Kʌrewari�K��rohtak�Ksirsa�Kƌsonipat�KŌyamunanagar�Kیbilaspur�K֌chamba�Kٌhamirpur�KՌkangra�K،kinnaur�Kӌkullu�KҌlahaul spiti�K׌mandi�KЌshimla�KԌsirmaur�Kьsolan�Kڌuna�K��anantnag�Kߌ	bandipore�K�	baramulla�K�budgam�K�doda�K�	ganderbal�K�jammu�K�kathua�K�kishtwar�K݌kulgam�K�kupwara�K�poonch�K�pulwama�K�rajouri�K�ramban�K�reasi�K�samba�Kތshopian�K܌srinagar�K�udhampur�K�bokaro�K��chatra�K��deoghar�M�dhanbad�M�dumka�K��east singhbhum�K�garhwa�M �giridih�M�godda�K��gumla�K��
hazaribagh�M�jamtara�K��khunti�K�koderma�K�latehar�K��	lohardaga�M�pakur�K��palamu�K��ramgarh�K��ranchi�M�	sahebganj�K��seraikela kharsawan�K��simdega�M�west singhbhum�M�bagalkot�M�bangalore rural�M	�bangalore urban�M&�bbmp�M�belgaum�M�bellary�M�bidar�M�chamarajanagar�M�chikamagalur�M#�chikkaballapur�M�chitradurga�M�dakshina kannada�M�
davanagere�M�dharwad�M�gadag�M�gulbarga�M!�hassan�M�haveri�M�kodagu�M�kolar�M�koppal�M"�mandya�M
�mysore�M�raichur�M$�
ramanagara�M�shimoga�M �tumkur�M�udupi�M�uttar kannada�M%�
vijayapura�M�yadgir�M-�	alappuzha�M3�	ernakulam�M2�idukki�M)�kannur�M'�	kasaragod�M*�kollam�M0�kottayam�M1�	kozhikode�M.�
malappuram�M4�palakkad�M,�pathanamthitta�M(�thiruvananthapuram�M/�thrissur�M+�wayanad�M5�kargil�M6�leh�M�agatti island�M7�lakshadweep�M@�agar�Me�	alirajpur�MN�anuppur�Mb�
ashoknagar�MR�balaghat�MW�barwani�Mj�betul�M_�bhind�M8�bhopal�MV�	burhanpur�MH�
chhatarpur�MQ�
chhindwara�MG�damoh�M^�datia�MD�dewas�MU�dhar�MP�dindori�M\�guna�M9�gwalior�Mi�harda�Mh�hoshangabad�M:�indore�M;�jabalpur�MT�jhabua�Ma�katni�MS�khandwa�MX�khargone�MO�mandla�M?�mandsaur�M[�morena�M`�narsinghpur�MC�neemuch�MF�panna�Mg�raisen�Mf�rajgarh�MB�ratlam�M<�rewa�M=�sagar�MM�satna�Md�sehore�M]�seoni�ML�shahdol�MA�shajapur�MZ�sheopur�MY�shivpuri�MK�sidhi�MJ�	singrauli�ME�	tikamgarh�M>�ujjain�MI�umaria�Mc�vidisha�M��
ahmednagar�Ml�akola�Mn�amravati�M��aurangabad �M��beed�Mr�bhandara�Mo�buldhana�M|�
chandrapur�M��dhule�M{�
gadchiroli�Mz�gondia�M��hingoli�M��jalgaon�M��jalna�Ms�kolhapur�M�latur�M��mumbai�Mm�nagpur�M~�nanded�M��	nandurbar�M��nashik�M}�	osmanabad�M��palghar�M��parbhani�Mk�pune�M��raigad�Mt�	ratnagiri�Mu�sangli�Mx�satara�Mv�
sindhudurg�Mw�solapur�M��thane�My�wardha�Mq�washim�Mp�yavatmal�M��	bishnupur�M��chandel�M��churachandpur�M��imphal east�M��imphal west�M��jiribam�M��kakching�M��kamjong�M��	kangpokpi�M��noney�M��pherzawl�M��senapati�M��
tamenglong�M��
tengnoupal�M��thoubal�M��ukhrul�M��east garo hills�M��east jaintia hills�M��east khasi hills�M��north garo hills�M��ri-bhoi�M��south garo hills�M��south west garo hills�M��south west khasi hills�M��west garo hills�M��west jaintia hills�M��west khasi hills�M��aizawl east�M��aizawl west�M��champhai�M��kolasib�M��	lawngtlai�M��lunglei�M��mamit�M��serchhip�M��siaha�M��dimapur�M��kiphire�M��kohima�M��longleng�M��
mokokchung�M��mon�M��peren�M��phek�M��tuensang�M��wokha�M��	zunheboto�M��angul�M��balangir�M��balasore�M��bargarh�M��bhadrak�M��boudh�M��cuttack�M��deogarh�M��	dhenkanal�M��gajapati�M��ganjam�M��jagatsinghpur�M��jajpur�M��
jharsuguda�M��	kalahandi�M��	kandhamal�M��
kendrapara�M��	kendujhar�M��khurda�M��koraput�M��
malkangiri�M��
mayurbhanj�M��nabarangpur�M��nayagarh�M��nuapada�M��puri�M��rayagada�M��	sambalpur�M��
subarnapur�M��
sundargarh�M��karaikal�M��mahe�M��
puducherry�M��yanam�M��amritsar�M��barnala�M��bathinda�M��faridkot�M��fatehgarh sahib�M��fazilka�M��ferozpur�M��	gurdaspur�M��
hoshiarpur�M��	jalandhar�M��
kapurthala�M��ludhiana�M��mansa�M��moga�M��	pathankot�M��patiala�M��	rup nagar�M��sangrur�M��	sas nagar�M��	sbs nagar�M��sri muktsar sahib�M��
tarn taran�M��ajmer�M �alwar�M�banswara�M�baran�M�barmer�M��	bharatpur�M�bhilwara�M��bikaner�M�bundi�M	�chittorgarh�M�churu�M��dausa�M�dholpur�M�	dungarpur�M�hanumangarh�M��jaipur i�M��	jaipur ii�M�	jaisalmer�M�jalore�M�jhalawar�M��	jhunjhunu�M��jodhpur�M�karauli�M��kota�M�nagaur�M�pali�M
�
pratapgarh�M�	rajsamand�M�sawai madhopur�M�sikar�M�sirohi�M��sri ganganagar�M�tonk�M��udaipur�M�east sikkim�M�north sikkim�M�south sikkim�M�west sikkim�M�
aranthangi�M+�ariyalur�MB�attur�M5�
chengalpet�M;�chennai�M
�cheyyar�M�
coimbatore�M#�	cuddalore�M6�
dharmapuri�M,�dindigul�M3�erode�M(�kallakurichi�M-�kanchipuram�M �kanyakumari�M/�karur�M�
kovilpatti�M2�krishnagiri�M�madurai�M@�nagapattinam�M.�namakkal�MA�nilgiris�M4�palani�M=�
paramakudi�M:�
perambalur�M?�poonamallee�M"�pudukkottai�M7�ramanathapuram�M�ranipet�M!�salem�M1�	sivaganga�MD�sivakasi�M'�tenkasi�M�	thanjavur�M9�theni�M*�thoothukudi (tuticorin)�M0�tiruchirappalli�M$�tirunelveli�M&�
tirupattur�M8�tiruppur�M<�
tiruvallur�M)�tiruvannamalai�M>�	tiruvarur�M�vellore�M�
viluppuram�M%�virudhunagar�MF�adilabad�MG�bhadradri kothagudem�ME�	hyderabad�MH�jagtial�MI�jangaon�MJ�jayashankar bhupalpally�MK�jogulamba gadwal�ML�	kamareddy�MM�
karimnagar�MN�khammam�MO�kumuram bheem�MP�mahabubabad�MQ�mahabubnagar�MR�
mancherial�MS�medak�MT�medchal�Md�mulugu�MU�nagarkurnool�MV�nalgonda�Me�
narayanpet�MW�nirmal�MX�	nizamabad�MY�
peddapalli�MZ�rajanna sircilla�M[�
rangareddy�M\�
sangareddy�M]�siddipet�M^�suryapet�M_�	vikarabad�M`�
wanaparthy�Ma�warangal(rural)�Mb�warangal(urban)�Mc�yadadri bhuvanagiri�Mf�dhalai�Mg�gomati�Mh�khowai�Mi�north tripura�Mj�
sepahijala�Mk�south tripura�Ml�unakoti�Mm�west tripura�Mn�agra�Mo�aligarh�Mq�ambedkar nagar�Mr�amethi�Ms�amroha�Mt�auraiya�M��ayodhya�Mu�azamgarh�Mv�badaun�Mw�baghpat�Mx�bahraich�My�
balarampur�Mz�ballia�M{�banda�M|�	barabanki�M}�bareilly�M~�basti�M��bhadohi�M�bijnour�M��bulandshahr�M��	chandauli�M��
chitrakoot�M��deoria�M��etah�M��etawah�M��farrukhabad�M��fatehpur�M��	firozabad�M��gautam buddha nagar�M��	ghaziabad�M��ghazipur�M��gonda�M��	gorakhpur�M��hamirpur�M��hapur�M��hardoi�M��hathras�M��jalaun�M��jaunpur�M��jhansi�M��kannauj�M��kanpur dehat�M��kanpur nagar�M��kasganj�M��	kaushambi�M��
kushinagar�M��lakhimpur kheri�M��lalitpur�M��lucknow�M��maharajganj�M��mahoba�M��mainpuri�M��mathura�M��mau�M��meerut�M��mirzapur�M��	moradabad�M��muzaffarnagar�M��pilibhit�M��
pratapgarh�Mp�	prayagraj�M��	raebareli�M��rampur�M��
saharanpur�M��sambhal�M��sant kabir nagar�M��shahjahanpur�M��shamli�M��	shravasti�M��siddharthnagar�M��sitapur�M��	sonbhadra�M��	sultanpur�M��unnao�M��varanasi�M��almora�M��	bageshwar�M��chamoli�M��	champawat�M��dehradun�M��haridwar�M��nainital�M��pauri garhwal�M��pithoragarh�M��rudraprayag�M��tehri garhwal�M��udham singh nagar�M��
uttarkashi�M��alipurduar district�M��bankura�M��basirhat hd (north 24 parganas)�M��birbhum�M��bishnupur hd (bankura)�M��cooch behar�M�
coochbehar�M��dakshin dinajpur�M��
darjeeling�M��!diamond harbor hd (s 24 parganas)�M��east bardhaman�M��hoogly�M��howrah�M��
jalpaiguri�M��jhargram�M��	kalimpong�M��kolkata�M��malda�M��murshidabad�M��nadia�M��nandigram hd (east medinipore)�M��north 24 parganas�M��paschim medinipore�M��purba medinipore�M��purulia�M��rampurhat hd (birbhum)�M��south 24 parganas�M��uttar dinajpur�M��west bardhaman�u.