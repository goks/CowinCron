���+      }�(K}�(�nicobar�K�north and middle andaman�K�south andaman�KuK}�(�	anantapur�K	�chittoor�K
�east godavari�K�guntur�K�krishna�K�kurnool�K�prakasam�K�sri potti sriramulu nellore�K�
srikakulam�K�visakhapatnam�K�vizianagaram�K�west godavari�K�ysr district, kadapa (cuddapah)�KuK}�(�anjaw�K�	changlang�K�dibang valley�K�east kameng�K�
east siang�K*�itanagar capital complex�K�kamle�K�	kra daadi�K�kurung kumey�K�	lepa rada�K!�lohit�K�longding�K(�lower dibang valley�K�lower siang�K�lower subansiri�K �namsai�K$�pakke kessang�K�
papum pare�K'�shi yomi�K#�siang�K%�tawang�K�tirap�K�upper siang�K"�upper subansiri�K)�west kameng�K�
west siang�K&uK}�(�baksa�K.�barpeta�K/�	biswanath�M��
bongaigaon�K9�cachar�KB�	charaideo�M��chirang�K:�darrang�K0�dhemaji�K>�dhubri�K;�	dibrugarh�K+�
dima hasao�KC�goalpara�K<�golaghat�K5�
hailakandi�KD�hojai�M��jorhat�K6�kamrup metropolitan�K1�kamrup rural�K2�karbi-anglong�K3�	karimganj�KE�	kokrajhar�K=�	lakhimpur�K?�majuli�M��morigaon�K7�nagaon�K8�nalbari�K4�	sivasagar�K,�sonitpur�K@�south salmara mankachar�M �tinsukia�K-�udalguri�KA�west karbi anglong�MuK}�(�araria�KJ�arwal�KN�
aurangabad�KM�banka�KS�	begusarai�Kb�	bhagalpur�KR�bhojpur�Kc�buxar�Kd�	darbhanga�K^�east champaran�Ki�gaya�KO�	gopalganj�Kh�jamui�Kk�	jehanabad�K[�kaimur�KP�katihar�KK�khagaria�Ke�
kishanganj�KL�
lakhisarai�KT�	madhepura�KF�	madhubani�K_�munger�KU�muzaffarpur�KV�nalanda�KZ�nawada�K\�patna�Ka�purnia�KI�rohtas�KQ�saharsa�KG�
samastipur�K`�saran�Kf�
sheikhpura�K]�sheohar�KW�	sitamarhi�KX�siwan�Kg�supaul�KH�vaishali�KY�west champaran�KjuK}��
chandigarh�KlsK}�(�balod�Kn�baloda bazar�Ko�	balrampur�Kp�bastar�Kq�bemetara�Kr�bijapur�Ks�bilaspur�Kt�	dantewada�Ku�dhamtari�Kv�durg�Kw�	gariaband�Kx�gaurela pendra marwahi �K��janjgir-champa�Ky�jashpur�Kz�kanker�K{�kawardha�K��	kondagaon�K|�korba�K}�koriya�K~�
mahasamund�K�mungeli�K��
narayanpur�K��raigarh�K��raipur�Km�rajnandgaon�K��sukma�K��surajpur�K��surguja�K�uK}��dadra and nagar haveli�K�sK%}�(�daman�K��diu�K�uK	}�(�central delhi�K��
east delhi�K��	new delhi�K��north delhi�K��north east delhi�K��north west delhi�K��shahdara�K��south delhi�K��south east delhi�K��south west delhi�K��
west delhi�K�uK
}�(�	north goa�K��	south goa�K�uK}�(�	ahmedabad�K��ahmedabad corporation�M�amreli�K��anand�K��aravalli�K��banaskantha�K��bharuch�K��	bhavnagar�K��bhavnagar corporation�M�botad�K��chhotaudepur�K��dahod�K��dang�K��devbhumi dwaraka�K��gandhinagar�K��gandhinagar corporation�M�gir somnath�K��jamnagar�K��jamnagar corporation�M�junagadh�K��junagadh corporation�M�kheda�K��kutch�K��	mahisagar�K��mehsana�K��morbi�K��narmada�K��navsari�K��
panchmahal�K��patan�K��	porbandar�K��rajkot�K��rajkot corporation�M�sabarkantha�K��surat�K��surat corporation�M�surendranagar�K��tapi�K��vadodara�K��vadodara corporation�M	�valsad�K�uK}�(�ambala�K��bhiwani�KȌcharkhi dadri�KɌ	faridabad�Kǌ	fatehabad�KČgurgaon�K��hisar�K��jhajjar�K��jind�Ǩkaithal�K��karnal�Kˌkurukshetra�K��mahendragarh�KΌnuh�K͌palwal�Kό	panchkula�K��panipat�KÌrewari�Kʌrohtak�K��sirsa�Ksonipat�Kƌyamunanagar�K�uK}�(�bilaspur�Kیchamba�K֌hamirpur�Kٌkangra�KՌkinnaur�K،kullu�Kӌlahaul spiti�KҌmandi�K׌shimla�KЌsirmaur�KԌsolan�Kьuna�K�uK}�(�anantnag�K��	bandipore�Kߌ	baramulla�K�budgam�K�doda�K�	ganderbal�K�jammu�K�kathua�K�kishtwar�K�kulgam�K݌kupwara�K�poonch�K�pulwama�K�rajouri�K�ramban�K�reasi�K�samba�K�shopian�Kތsrinagar�K܌udhampur�K�uK}�(�bokaro�K�chatra�K��deoghar�K��dhanbad�M�dumka�M�east singhbhum�K��garhwa�K�giridih�M �godda�M�gumla�K��
hazaribagh�K��jamtara�M�khunti�K��koderma�K�latehar�K�	lohardaga�K��pakur�M�palamu�K��ramgarh�K��ranchi�K��	sahebganj�M�seraikela kharsawan�K��simdega�K��west singhbhum�MuK}�(�bagalkot�M�bangalore rural�M�bangalore urban�M	�bbmp�M&�belgaum�M�bellary�M�bidar�M�chamarajanagar�M�chikamagalur�M�chikkaballapur�M#�chitradurga�M�dakshina kannada�M�
davanagere�M�dharwad�M�gadag�M�gulbarga�M�hassan�M!�haveri�M�kodagu�M�kolar�M�koppal�M�mandya�M"�mysore�M
�raichur�M�
ramanagara�M$�shimoga�M�tumkur�M �udupi�M�uttar kannada�M�
vijayapura�M%�yadgir�MuK}�(�	alappuzha�M-�	ernakulam�M3�idukki�M2�kannur�M)�	kasaragod�M'�kollam�M*�kottayam�M0�	kozhikode�M1�
malappuram�M.�palakkad�M4�pathanamthitta�M,�thiruvananthapuram�M(�thrissur�M/�wayanad�M+uK}�(�kargil�M5�leh�M6uK}�(�agatti island�M�lakshadweep�M7uK}�(�agar�M@�	alirajpur�Me�anuppur�MN�
ashoknagar�Mb�balaghat�MR�barwani�MW�betul�Mj�bhind�M_�bhopal�M8�	burhanpur�MV�
chhatarpur�MH�
chhindwara�MQ�damoh�MG�datia�M^�dewas�MD�dhar�MU�dindori�MP�guna�M\�gwalior�M9�harda�Mi�hoshangabad�Mh�indore�M:�jabalpur�M;�jhabua�MT�katni�Ma�khandwa�MS�khargone�MX�mandla�MO�mandsaur�M?�morena�M[�narsinghpur�M`�neemuch�MC�panna�MF�raisen�Mg�rajgarh�Mf�ratlam�MB�rewa�M<�sagar�M=�satna�MM�sehore�Md�seoni�M]�shahdol�ML�shajapur�MA�sheopur�MZ�shivpuri�MY�sidhi�MK�	singrauli�MJ�	tikamgarh�ME�ujjain�M>�umaria�MI�vidisha�McuK}�(�
ahmednagar�M��akola�Ml�amravati�Mn�aurangabad �M��beed�M��bhandara�Mr�buldhana�Mo�
chandrapur�M|�dhule�M��
gadchiroli�M{�gondia�Mz�hingoli�M��jalgaon�M��jalna�M��kolhapur�Ms�latur�M�mumbai�M��nagpur�Mm�nanded�M~�	nandurbar�M��nashik�M��	osmanabad�M}�palghar�M��parbhani�M��pune�Mk�raigad�M��	ratnagiri�Mt�sangli�Mu�satara�Mx�
sindhudurg�Mv�solapur�Mw�thane�M��wardha�My�washim�Mq�yavatmal�MpuK}�(�	bishnupur�M��chandel�M��churachandpur�M��imphal east�M��imphal west�M��jiribam�M��kakching�M��kamjong�M��	kangpokpi�M��noney�M��pherzawl�M��senapati�M��
tamenglong�M��
tengnoupal�M��thoubal�M��ukhrul�M�uK}�(�east garo hills�M��east jaintia hills�M��east khasi hills�M��north garo hills�M��ri-bhoi�M��south garo hills�M��south west garo hills�M��south west khasi hills�M��west garo hills�M��west jaintia hills�M��west khasi hills�M�uK}�(�aizawl east�M��aizawl west�M��champhai�M��kolasib�M��	lawngtlai�M��lunglei�M��mamit�M��serchhip�M��siaha�M�uK}�(�dimapur�M��kiphire�M��kohima�M��longleng�M��
mokokchung�M��mon�M��peren�M��phek�M��tuensang�M��wokha�M��	zunheboto�M�uK}�(�angul�M��balangir�M��balasore�M��bargarh�M��bhadrak�M��boudh�M��cuttack�M��deogarh�M��	dhenkanal�M��gajapati�M��ganjam�M��jagatsinghpur�M��jajpur�M��
jharsuguda�M��	kalahandi�M��	kandhamal�M��
kendrapara�M��	kendujhar�M��khurda�M��koraput�M��
malkangiri�M��
mayurbhanj�M��nabarangpur�M��nayagarh�M��nuapada�M��puri�M��rayagada�M��	sambalpur�M��
subarnapur�M��
sundargarh�M�uK}�(�karaikal�M��mahe�M��
puducherry�M��yanam�M�uK}�(�amritsar�M��barnala�M��bathinda�M��faridkot�M��fatehgarh sahib�M��fazilka�M��ferozpur�M��	gurdaspur�M��
hoshiarpur�M��	jalandhar�M��
kapurthala�M��ludhiana�M��mansa�M��moga�M��	pathankot�M��patiala�M��	rup nagar�M��sangrur�M��	sas nagar�M��	sbs nagar�M��sri muktsar sahib�M��
tarn taran�M�uK}�(�ajmer�M��alwar�M �banswara�M�baran�M�barmer�M�	bharatpur�M��bhilwara�M�bikaner�M��bundi�M�chittorgarh�M	�churu�M�dausa�M��dholpur�M�	dungarpur�M�hanumangarh�M�jaipur i�M��	jaipur ii�M��	jaisalmer�M�jalore�M�jhalawar�M�	jhunjhunu�M��jodhpur�M��karauli�M�kota�M��nagaur�M�pali�M�
pratapgarh�M
�	rajsamand�M�sawai madhopur�M�sikar�M�sirohi�M�sri ganganagar�M��tonk�M�udaipur�M�uK}�(�east sikkim�M�north sikkim�M�south sikkim�M�west sikkim�MuK}�(�
aranthangi�M�ariyalur�M+�attur�MB�
chengalpet�M5�chennai�M;�cheyyar�M
�
coimbatore�M�	cuddalore�M#�
dharmapuri�M6�dindigul�M,�erode�M3�kallakurichi�M(�kanchipuram�M-�kanyakumari�M �karur�M/�
kovilpatti�M�krishnagiri�M2�madurai�M�nagapattinam�M@�namakkal�M.�nilgiris�MA�palani�M4�
paramakudi�M=�
perambalur�M:�poonamallee�M?�pudukkottai�M"�ramanathapuram�M7�ranipet�M�salem�M!�	sivaganga�M1�sivakasi�MD�tenkasi�M'�	thanjavur�M�theni�M9�thoothukudi (tuticorin)�M*�tiruchirappalli�M0�tirunelveli�M$�
tirupattur�M&�tiruppur�M8�
tiruvallur�M<�tiruvannamalai�M)�	tiruvarur�M>�vellore�M�
viluppuram�M�virudhunagar�M%uK }�(�adilabad�MF�bhadradri kothagudem�MG�	hyderabad�ME�jagtial�MH�jangaon�MI�jayashankar bhupalpally�MJ�jogulamba gadwal�MK�	kamareddy�ML�
karimnagar�MM�khammam�MN�kumuram bheem�MO�mahabubabad�MP�mahabubnagar�MQ�
mancherial�MR�medak�MS�medchal�MT�mulugu�Md�nagarkurnool�MU�nalgonda�MV�
narayanpet�Me�nirmal�MW�	nizamabad�MX�
peddapalli�MY�rajanna sircilla�MZ�
rangareddy�M[�
sangareddy�M\�siddipet�M]�suryapet�M^�	vikarabad�M_�
wanaparthy�M`�warangal(rural)�Ma�warangal(urban)�Mb�yadadri bhuvanagiri�McuK!}�(�dhalai�Mf�gomati�Mg�khowai�Mh�north tripura�Mi�
sepahijala�Mj�south tripura�Mk�unakoti�Ml�west tripura�MmuK"}�(�agra�Mn�aligarh�Mo�ambedkar nagar�Mq�amethi�Mr�amroha�Ms�auraiya�Mt�ayodhya�M��azamgarh�Mu�badaun�Mv�baghpat�Mw�bahraich�Mx�
balarampur�My�ballia�Mz�banda�M{�	barabanki�M|�bareilly�M}�basti�M~�bhadohi�M��bijnour�M�bulandshahr�M��	chandauli�M��
chitrakoot�M��deoria�M��etah�M��etawah�M��farrukhabad�M��fatehpur�M��	firozabad�M��gautam buddha nagar�M��	ghaziabad�M��ghazipur�M��gonda�M��	gorakhpur�M��hamirpur�M��hapur�M��hardoi�M��hathras�M��jalaun�M��jaunpur�M��jhansi�M��kannauj�M��kanpur dehat�M��kanpur nagar�M��kasganj�M��	kaushambi�M��
kushinagar�M��lakhimpur kheri�M��lalitpur�M��lucknow�M��maharajganj�M��mahoba�M��mainpuri�M��mathura�M��mau�M��meerut�M��mirzapur�M��	moradabad�M��muzaffarnagar�M��pilibhit�M��
pratapgarh�M��	prayagraj�Mp�	raebareli�M��rampur�M��
saharanpur�M��sambhal�M��sant kabir nagar�M��shahjahanpur�M��shamli�M��	shravasti�M��siddharthnagar�M��sitapur�M��	sonbhadra�M��	sultanpur�M��unnao�M��varanasi�M�uK#}�(�almora�M��	bageshwar�M��chamoli�M��	champawat�M��dehradun�M��haridwar�M��nainital�M��pauri garhwal�M��pithoragarh�M��rudraprayag�M��tehri garhwal�M��udham singh nagar�M��
uttarkashi�M�uK$}�(�alipurduar district�M��bankura�M��basirhat hd (north 24 parganas)�M��birbhum�M��bishnupur hd (bankura)�M��cooch behar�M��
coochbehar�M�dakshin dinajpur�M��
darjeeling�M��!diamond harbor hd (s 24 parganas)�M��east bardhaman�M��hoogly�M��howrah�M��
jalpaiguri�M��jhargram�M��	kalimpong�M��kolkata�M��malda�M��murshidabad�M��nadia�M��nandigram hd (east medinipore)�M��north 24 parganas�M��paschim medinipore�M��purba medinipore�M��purulia�M��rampurhat hd (birbhum)�M��south 24 parganas�M��uttar dinajpur�M��west bardhaman�M�uu.